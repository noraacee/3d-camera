// nios_system.v

// Generated using ACDS version 13.0sp1 232 at 2015.04.08.21:18:30

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clock_50_clk,                //       clock_50.clk
		input  wire        reset_50_reset_n,            //       reset_50.reset_n
		input  wire        video_decoder_TD_CLK27,      //  video_decoder.TD_CLK27
		input  wire [7:0]  video_decoder_TD_DATA,       //               .TD_DATA
		input  wire        video_decoder_TD_HS,         //               .TD_HS
		input  wire        video_decoder_TD_VS,         //               .TD_VS
		input  wire        video_decoder_clk27_reset,   //               .clk27_reset
		output wire        video_decoder_TD_RESET,      //               .TD_RESET
		output wire        video_decoder_overflow_flag, //               .overflow_flag
		inout  wire [15:0] sram_DQ,                     //           sram.DQ
		output wire [17:0] sram_ADDR,                   //               .ADDR
		output wire        sram_LB_N,                   //               .LB_N
		output wire        sram_UB_N,                   //               .UB_N
		output wire        sram_CE_N,                   //               .CE_N
		output wire        sram_OE_N,                   //               .OE_N
		output wire        sram_WE_N,                   //               .WE_N
		output wire        vga_controller_CLK,          // vga_controller.CLK
		output wire        vga_controller_HS,           //               .HS
		output wire        vga_controller_VS,           //               .VS
		output wire        vga_controller_BLANK,        //               .BLANK
		output wire        vga_controller_SYNC,         //               .SYNC
		output wire [9:0]  vga_controller_R,            //               .R
		output wire [9:0]  vga_controller_G,            //               .G
		output wire [9:0]  vga_controller_B,            //               .B
		output wire        threedlizer_reset_out,       //    threedlizer.reset_out
		input  wire        threedlizer_pixel_r_ready,   //               .pixel_r_ready
		input  wire [4:0]  threedlizer_pixel_r,         //               .pixel_r
		input  wire [17:0] threedlizer_pixel_offset,    //               .pixel_offset
		output wire        threedlizer_pixel_r_done,    //               .pixel_r_done
		output wire [17:0] threedlizer_red_led,         //               .red_led
		input  wire        threedlizer_clk_in,          //               .clk_in
		input  wire        buffer_reader_clk_in,        //  buffer_reader.clk_in
		input  wire        buffer_reader_pixel_set,     //               .pixel_set
		input  wire [17:0] buffer_reader_pixel_offset,  //               .pixel_offset
		output wire        buffer_reader_pixel_ready,   //               .pixel_ready
		output wire [15:0] buffer_reader_pixel,         //               .pixel
		output wire [1:0]  buffer_reader_red_led        //               .red_led
	);

	wire         clocks_sys_clk_clk;                                                                               // clocks:sys_clk -> [3Dlizer:clk, 3Dlizer_avalon_master_r_translator:clk, 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:clk, 3Dlizer_avalon_master_w_translator:clk, 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, buffer_reader:clk, buffer_reader_avalon_master_translator:clk, buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:clk, chroma_resampler:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_mux:clk, color_space_converter:clk, dual_clock_fifo:clk_stream_in, id_router:clk, p_buffer:clk, p_buffer_avalon_sram_slave_translator:clk, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, p_buffer_dma:clk, p_buffer_dma_avalon_pixel_dma_master_translator:clk, p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, p_rgb_resampler:clk, p_scaler:clk, rsp_xbar_demux:clk, rst_controller_001:clk, v_clipper:clk, v_decoder:clk, v_dma_controller:clk, v_dma_controller_avalon_dma_master_translator:clk, v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, v_rgb_resampler:clk, v_scaler:clk]
	wire         v_decoder_avalon_decoder_source_endofpacket;                                                      // v_decoder:stream_out_endofpacket -> chroma_resampler:stream_in_endofpacket
	wire         v_decoder_avalon_decoder_source_valid;                                                            // v_decoder:stream_out_valid -> chroma_resampler:stream_in_valid
	wire         v_decoder_avalon_decoder_source_startofpacket;                                                    // v_decoder:stream_out_startofpacket -> chroma_resampler:stream_in_startofpacket
	wire  [15:0] v_decoder_avalon_decoder_source_data;                                                             // v_decoder:stream_out_data -> chroma_resampler:stream_in_data
	wire         v_decoder_avalon_decoder_source_ready;                                                            // chroma_resampler:stream_in_ready -> v_decoder:stream_out_ready
	wire         chroma_resampler_avalon_chroma_source_endofpacket;                                                // chroma_resampler:stream_out_endofpacket -> color_space_converter:stream_in_endofpacket
	wire         chroma_resampler_avalon_chroma_source_valid;                                                      // chroma_resampler:stream_out_valid -> color_space_converter:stream_in_valid
	wire         chroma_resampler_avalon_chroma_source_startofpacket;                                              // chroma_resampler:stream_out_startofpacket -> color_space_converter:stream_in_startofpacket
	wire  [23:0] chroma_resampler_avalon_chroma_source_data;                                                       // chroma_resampler:stream_out_data -> color_space_converter:stream_in_data
	wire         chroma_resampler_avalon_chroma_source_ready;                                                      // color_space_converter:stream_in_ready -> chroma_resampler:stream_out_ready
	wire         color_space_converter_avalon_csc_source_endofpacket;                                              // color_space_converter:stream_out_endofpacket -> v_rgb_resampler:stream_in_endofpacket
	wire         color_space_converter_avalon_csc_source_valid;                                                    // color_space_converter:stream_out_valid -> v_rgb_resampler:stream_in_valid
	wire         color_space_converter_avalon_csc_source_startofpacket;                                            // color_space_converter:stream_out_startofpacket -> v_rgb_resampler:stream_in_startofpacket
	wire  [23:0] color_space_converter_avalon_csc_source_data;                                                     // color_space_converter:stream_out_data -> v_rgb_resampler:stream_in_data
	wire         color_space_converter_avalon_csc_source_ready;                                                    // v_rgb_resampler:stream_in_ready -> color_space_converter:stream_out_ready
	wire         v_rgb_resampler_avalon_rgb_source_endofpacket;                                                    // v_rgb_resampler:stream_out_endofpacket -> v_clipper:stream_in_endofpacket
	wire         v_rgb_resampler_avalon_rgb_source_valid;                                                          // v_rgb_resampler:stream_out_valid -> v_clipper:stream_in_valid
	wire         v_rgb_resampler_avalon_rgb_source_startofpacket;                                                  // v_rgb_resampler:stream_out_startofpacket -> v_clipper:stream_in_startofpacket
	wire  [15:0] v_rgb_resampler_avalon_rgb_source_data;                                                           // v_rgb_resampler:stream_out_data -> v_clipper:stream_in_data
	wire         v_rgb_resampler_avalon_rgb_source_ready;                                                          // v_clipper:stream_in_ready -> v_rgb_resampler:stream_out_ready
	wire         v_clipper_avalon_clipper_source_endofpacket;                                                      // v_clipper:stream_out_endofpacket -> v_scaler:stream_in_endofpacket
	wire         v_clipper_avalon_clipper_source_valid;                                                            // v_clipper:stream_out_valid -> v_scaler:stream_in_valid
	wire         v_clipper_avalon_clipper_source_startofpacket;                                                    // v_clipper:stream_out_startofpacket -> v_scaler:stream_in_startofpacket
	wire  [15:0] v_clipper_avalon_clipper_source_data;                                                             // v_clipper:stream_out_data -> v_scaler:stream_in_data
	wire         v_clipper_avalon_clipper_source_ready;                                                            // v_scaler:stream_in_ready -> v_clipper:stream_out_ready
	wire         v_scaler_avalon_scaler_source_endofpacket;                                                        // v_scaler:stream_out_endofpacket -> v_dma_controller:stream_endofpacket
	wire         v_scaler_avalon_scaler_source_valid;                                                              // v_scaler:stream_out_valid -> v_dma_controller:stream_valid
	wire         v_scaler_avalon_scaler_source_startofpacket;                                                      // v_scaler:stream_out_startofpacket -> v_dma_controller:stream_startofpacket
	wire  [15:0] v_scaler_avalon_scaler_source_data;                                                               // v_scaler:stream_out_data -> v_dma_controller:stream_data
	wire         v_scaler_avalon_scaler_source_ready;                                                              // v_dma_controller:stream_ready -> v_scaler:stream_out_ready
	wire         p_buffer_dma_avalon_pixel_source_endofpacket;                                                     // p_buffer_dma:stream_endofpacket -> p_rgb_resampler:stream_in_endofpacket
	wire         p_buffer_dma_avalon_pixel_source_valid;                                                           // p_buffer_dma:stream_valid -> p_rgb_resampler:stream_in_valid
	wire         p_buffer_dma_avalon_pixel_source_startofpacket;                                                   // p_buffer_dma:stream_startofpacket -> p_rgb_resampler:stream_in_startofpacket
	wire  [15:0] p_buffer_dma_avalon_pixel_source_data;                                                            // p_buffer_dma:stream_data -> p_rgb_resampler:stream_in_data
	wire         p_buffer_dma_avalon_pixel_source_ready;                                                           // p_rgb_resampler:stream_in_ready -> p_buffer_dma:stream_ready
	wire         p_rgb_resampler_avalon_rgb_source_endofpacket;                                                    // p_rgb_resampler:stream_out_endofpacket -> p_scaler:stream_in_endofpacket
	wire         p_rgb_resampler_avalon_rgb_source_valid;                                                          // p_rgb_resampler:stream_out_valid -> p_scaler:stream_in_valid
	wire         p_rgb_resampler_avalon_rgb_source_startofpacket;                                                  // p_rgb_resampler:stream_out_startofpacket -> p_scaler:stream_in_startofpacket
	wire  [29:0] p_rgb_resampler_avalon_rgb_source_data;                                                           // p_rgb_resampler:stream_out_data -> p_scaler:stream_in_data
	wire         p_rgb_resampler_avalon_rgb_source_ready;                                                          // p_scaler:stream_in_ready -> p_rgb_resampler:stream_out_ready
	wire         clocks_vga_clk_clk;                                                                               // clocks:VGA_CLK -> [dual_clock_fifo:clk_stream_out, rst_controller_002:clk, vga_controller:clk]
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                              // dual_clock_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                                                    // dual_clock_fifo:stream_out_valid -> vga_controller:valid
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                            // dual_clock_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                                                     // dual_clock_fifo:stream_out_data -> vga_controller:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                                                    // vga_controller:ready -> dual_clock_fifo:stream_out_ready
	wire         p_scaler_avalon_scaler_source_endofpacket;                                                        // p_scaler:stream_out_endofpacket -> dual_clock_fifo:stream_in_endofpacket
	wire         p_scaler_avalon_scaler_source_valid;                                                              // p_scaler:stream_out_valid -> dual_clock_fifo:stream_in_valid
	wire         p_scaler_avalon_scaler_source_startofpacket;                                                      // p_scaler:stream_out_startofpacket -> dual_clock_fifo:stream_in_startofpacket
	wire  [29:0] p_scaler_avalon_scaler_source_data;                                                               // p_scaler:stream_out_data -> dual_clock_fifo:stream_in_data
	wire         p_scaler_avalon_scaler_source_ready;                                                              // dual_clock_fifo:stream_in_ready -> p_scaler:stream_out_ready
	wire         p_buffer_dma_avalon_pixel_dma_master_waitrequest;                                                 // p_buffer_dma_avalon_pixel_dma_master_translator:av_waitrequest -> p_buffer_dma:master_waitrequest
	wire  [31:0] p_buffer_dma_avalon_pixel_dma_master_address;                                                     // p_buffer_dma:master_address -> p_buffer_dma_avalon_pixel_dma_master_translator:av_address
	wire         p_buffer_dma_avalon_pixel_dma_master_lock;                                                        // p_buffer_dma:master_arbiterlock -> p_buffer_dma_avalon_pixel_dma_master_translator:av_lock
	wire         p_buffer_dma_avalon_pixel_dma_master_read;                                                        // p_buffer_dma:master_read -> p_buffer_dma_avalon_pixel_dma_master_translator:av_read
	wire  [15:0] p_buffer_dma_avalon_pixel_dma_master_readdata;                                                    // p_buffer_dma_avalon_pixel_dma_master_translator:av_readdata -> p_buffer_dma:master_readdata
	wire         p_buffer_dma_avalon_pixel_dma_master_readdatavalid;                                               // p_buffer_dma_avalon_pixel_dma_master_translator:av_readdatavalid -> p_buffer_dma:master_readdatavalid
	wire         v_dma_controller_avalon_dma_master_waitrequest;                                                   // v_dma_controller_avalon_dma_master_translator:av_waitrequest -> v_dma_controller:master_waitrequest
	wire  [15:0] v_dma_controller_avalon_dma_master_writedata;                                                     // v_dma_controller:master_writedata -> v_dma_controller_avalon_dma_master_translator:av_writedata
	wire  [31:0] v_dma_controller_avalon_dma_master_address;                                                       // v_dma_controller:master_address -> v_dma_controller_avalon_dma_master_translator:av_address
	wire         v_dma_controller_avalon_dma_master_write;                                                         // v_dma_controller:master_write -> v_dma_controller_avalon_dma_master_translator:av_write
	wire         id3dlizer_avalon_master_w_waitrequest;                                                            // 3Dlizer_avalon_master_w_translator:av_waitrequest -> 3Dlizer:master_w_wait
	wire  [31:0] id3dlizer_avalon_master_w_address;                                                                // 3Dlizer:master_w_addr -> 3Dlizer_avalon_master_w_translator:av_address
	wire  [15:0] id3dlizer_avalon_master_w_writedata;                                                              // 3Dlizer:master_wd -> 3Dlizer_avalon_master_w_translator:av_writedata
	wire         id3dlizer_avalon_master_w_write;                                                                  // 3Dlizer:master_wr_en -> 3Dlizer_avalon_master_w_translator:av_write
	wire   [1:0] id3dlizer_avalon_master_w_byteenable;                                                             // 3Dlizer:master_w_be -> 3Dlizer_avalon_master_w_translator:av_byteenable
	wire         id3dlizer_avalon_master_r_waitrequest;                                                            // 3Dlizer_avalon_master_r_translator:av_waitrequest -> 3Dlizer:master_r_wait
	wire  [31:0] id3dlizer_avalon_master_r_address;                                                                // 3Dlizer:master_r_addr -> 3Dlizer_avalon_master_r_translator:av_address
	wire         id3dlizer_avalon_master_r_read;                                                                   // 3Dlizer:master_rd_en -> 3Dlizer_avalon_master_r_translator:av_read
	wire  [15:0] id3dlizer_avalon_master_r_readdata;                                                               // 3Dlizer_avalon_master_r_translator:av_readdata -> 3Dlizer:master_rd
	wire   [1:0] id3dlizer_avalon_master_r_byteenable;                                                             // 3Dlizer:master_r_be -> 3Dlizer_avalon_master_r_translator:av_byteenable
	wire         buffer_reader_avalon_master_waitrequest;                                                          // buffer_reader_avalon_master_translator:av_waitrequest -> buffer_reader:master_r_wait
	wire  [31:0] buffer_reader_avalon_master_address;                                                              // buffer_reader:master_r_addr -> buffer_reader_avalon_master_translator:av_address
	wire         buffer_reader_avalon_master_read;                                                                 // buffer_reader:master_rd_en -> buffer_reader_avalon_master_translator:av_read
	wire  [15:0] buffer_reader_avalon_master_readdata;                                                             // buffer_reader_avalon_master_translator:av_readdata -> buffer_reader:master_rd
	wire   [1:0] buffer_reader_avalon_master_byteenable;                                                           // buffer_reader:master_r_be -> buffer_reader_avalon_master_translator:av_byteenable
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                              // p_buffer_avalon_sram_slave_translator:av_writedata -> p_buffer:writedata
	wire  [17:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                // p_buffer_avalon_sram_slave_translator:av_address -> p_buffer:address
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                  // p_buffer_avalon_sram_slave_translator:av_write -> p_buffer:write
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                   // p_buffer_avalon_sram_slave_translator:av_read -> p_buffer:read
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                               // p_buffer:readdata -> p_buffer_avalon_sram_slave_translator:av_readdata
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                          // p_buffer:readdatavalid -> p_buffer_avalon_sram_slave_translator:av_readdatavalid
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                             // p_buffer_avalon_sram_slave_translator:av_byteenable -> p_buffer:byteenable
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;            // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> p_buffer_dma_avalon_pixel_dma_master_translator:uav_waitrequest
	wire   [1:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;             // p_buffer_dma_avalon_pixel_dma_master_translator:uav_burstcount -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;              // p_buffer_dma_avalon_pixel_dma_master_translator:uav_writedata -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                // p_buffer_dma_avalon_pixel_dma_master_translator:uav_address -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                   // p_buffer_dma_avalon_pixel_dma_master_translator:uav_lock -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                  // p_buffer_dma_avalon_pixel_dma_master_translator:uav_write -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                   // p_buffer_dma_avalon_pixel_dma_master_translator:uav_read -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;               // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> p_buffer_dma_avalon_pixel_dma_master_translator:uav_readdata
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;            // p_buffer_dma_avalon_pixel_dma_master_translator:uav_debugaccess -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;             // p_buffer_dma_avalon_pixel_dma_master_translator:uav_byteenable -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;          // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> p_buffer_dma_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;              // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> v_dma_controller_avalon_dma_master_translator:uav_waitrequest
	wire   [1:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;               // v_dma_controller_avalon_dma_master_translator:uav_burstcount -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;                // v_dma_controller_avalon_dma_master_translator:uav_writedata -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                  // v_dma_controller_avalon_dma_master_translator:uav_address -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                     // v_dma_controller_avalon_dma_master_translator:uav_lock -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                    // v_dma_controller_avalon_dma_master_translator:uav_write -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                     // v_dma_controller_avalon_dma_master_translator:uav_read -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                 // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> v_dma_controller_avalon_dma_master_translator:uav_readdata
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;              // v_dma_controller_avalon_dma_master_translator:uav_debugaccess -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;               // v_dma_controller_avalon_dma_master_translator:uav_byteenable -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;            // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> v_dma_controller_avalon_dma_master_translator:uav_readdatavalid
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_waitrequest;                       // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_waitrequest -> 3Dlizer_avalon_master_w_translator:uav_waitrequest
	wire   [1:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_burstcount;                        // 3Dlizer_avalon_master_w_translator:uav_burstcount -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_writedata;                         // 3Dlizer_avalon_master_w_translator:uav_writedata -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_address;                           // 3Dlizer_avalon_master_w_translator:uav_address -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_address
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_lock;                              // 3Dlizer_avalon_master_w_translator:uav_lock -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_lock
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_write;                             // 3Dlizer_avalon_master_w_translator:uav_write -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_write
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_read;                              // 3Dlizer_avalon_master_w_translator:uav_read -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdata;                          // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_readdata -> 3Dlizer_avalon_master_w_translator:uav_readdata
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_debugaccess;                       // 3Dlizer_avalon_master_w_translator:uav_debugaccess -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_byteenable;                        // 3Dlizer_avalon_master_w_translator:uav_byteenable -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_byteenable
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdatavalid;                     // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:av_readdatavalid -> 3Dlizer_avalon_master_w_translator:uav_readdatavalid
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_waitrequest;                       // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_waitrequest -> 3Dlizer_avalon_master_r_translator:uav_waitrequest
	wire   [1:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_burstcount;                        // 3Dlizer_avalon_master_r_translator:uav_burstcount -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_writedata;                         // 3Dlizer_avalon_master_r_translator:uav_writedata -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_address;                           // 3Dlizer_avalon_master_r_translator:uav_address -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_address
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_lock;                              // 3Dlizer_avalon_master_r_translator:uav_lock -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_lock
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_write;                             // 3Dlizer_avalon_master_r_translator:uav_write -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_write
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_read;                              // 3Dlizer_avalon_master_r_translator:uav_read -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdata;                          // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_readdata -> 3Dlizer_avalon_master_r_translator:uav_readdata
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_debugaccess;                       // 3Dlizer_avalon_master_r_translator:uav_debugaccess -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_byteenable;                        // 3Dlizer_avalon_master_r_translator:uav_byteenable -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_byteenable
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdatavalid;                     // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:av_readdatavalid -> 3Dlizer_avalon_master_r_translator:uav_readdatavalid
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_waitrequest;                     // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> buffer_reader_avalon_master_translator:uav_waitrequest
	wire   [1:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_burstcount;                      // buffer_reader_avalon_master_translator:uav_burstcount -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_writedata;                       // buffer_reader_avalon_master_translator:uav_writedata -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_address;                         // buffer_reader_avalon_master_translator:uav_address -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_lock;                            // buffer_reader_avalon_master_translator:uav_lock -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_write;                           // buffer_reader_avalon_master_translator:uav_write -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_read;                            // buffer_reader_avalon_master_translator:uav_read -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_readdata;                        // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> buffer_reader_avalon_master_translator:uav_readdata
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_debugaccess;                     // buffer_reader_avalon_master_translator:uav_debugaccess -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_byteenable;                      // buffer_reader_avalon_master_translator:uav_byteenable -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid;                   // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> buffer_reader_avalon_master_translator:uav_readdatavalid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // p_buffer_avalon_sram_slave_translator:uav_waitrequest -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> p_buffer_avalon_sram_slave_translator:uav_burstcount
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> p_buffer_avalon_sram_slave_translator:uav_writedata
	wire  [31:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> p_buffer_avalon_sram_slave_translator:uav_address
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> p_buffer_avalon_sram_slave_translator:uav_write
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> p_buffer_avalon_sram_slave_translator:uav_lock
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> p_buffer_avalon_sram_slave_translator:uav_read
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // p_buffer_avalon_sram_slave_translator:uav_readdata -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // p_buffer_avalon_sram_slave_translator:uav_readdatavalid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> p_buffer_avalon_sram_slave_translator:uav_debugaccess
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> p_buffer_avalon_sram_slave_translator:uav_byteenable
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [17:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;   // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;         // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket; // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [83:0] p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;          // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;         // addr_router:sink_ready -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;     // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;           // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;   // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [83:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;            // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;           // addr_router_001:sink_ready -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_endofpacket;              // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_valid;                    // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_startofpacket;            // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [83:0] id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_data;                     // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router_002:sink_ready -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:cp_ready
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket;              // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid;                    // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket;            // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [83:0] id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data;                     // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router_003:sink_ready -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:cp_ready
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;            // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                  // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;          // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [83:0] buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                   // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire         buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_004:sink_ready -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [83:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> clocks:reset
	wire         rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [3Dlizer:reset_in, 3Dlizer_avalon_master_r_translator:reset, 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:reset, 3Dlizer_avalon_master_w_translator:reset, 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, buffer_reader:rst, buffer_reader_avalon_master_translator:reset, buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:reset, chroma_resampler:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, color_space_converter:reset, dual_clock_fifo:reset_stream_in, id_router:reset, p_buffer:reset, p_buffer_avalon_sram_slave_translator:reset, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, p_buffer_dma:reset, p_buffer_dma_avalon_pixel_dma_master_translator:reset, p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, p_rgb_resampler:reset, p_scaler:reset, rsp_xbar_demux:reset, v_clipper:reset, v_decoder:reset, v_dma_controller:reset, v_dma_controller_avalon_dma_master_translator:reset, v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, v_rgb_resampler:reset, v_scaler:reset]
	wire         rst_controller_002_reset_out_reset;                                                               // rst_controller_002:reset_out -> [dual_clock_fifo:reset_stream_out, vga_controller:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [4:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [4:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux:sink2_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux:sink2_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux:sink2_startofpacket
	wire  [83:0] cmd_xbar_demux_002_src0_data;                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux:sink2_data
	wire   [4:0] cmd_xbar_demux_002_src0_channel;                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux:sink2_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                    // cmd_xbar_mux:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                              // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux:sink3_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                    // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux:sink3_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                            // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux:sink3_startofpacket
	wire  [83:0] cmd_xbar_demux_003_src0_data;                                                                     // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux:sink3_data
	wire   [4:0] cmd_xbar_demux_003_src0_channel;                                                                  // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux:sink3_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                    // cmd_xbar_mux:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire         cmd_xbar_demux_004_src0_endofpacket;                                                              // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux:sink4_endofpacket
	wire         cmd_xbar_demux_004_src0_valid;                                                                    // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux:sink4_valid
	wire         cmd_xbar_demux_004_src0_startofpacket;                                                            // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux:sink4_startofpacket
	wire  [83:0] cmd_xbar_demux_004_src0_data;                                                                     // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux:sink4_data
	wire   [4:0] cmd_xbar_demux_004_src0_channel;                                                                  // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux:sink4_channel
	wire         cmd_xbar_demux_004_src0_ready;                                                                    // cmd_xbar_mux:sink4_ready -> cmd_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src2_endofpacket;                                                                  // rsp_xbar_demux:src2_endofpacket -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src2_valid;                                                                        // rsp_xbar_demux:src2_valid -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src2_startofpacket;                                                                // rsp_xbar_demux:src2_startofpacket -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_demux_src2_data;                                                                         // rsp_xbar_demux:src2_data -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] rsp_xbar_demux_src2_channel;                                                                      // rsp_xbar_demux:src2_channel -> 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src3_endofpacket;                                                                  // rsp_xbar_demux:src3_endofpacket -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src3_valid;                                                                        // rsp_xbar_demux:src3_valid -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src3_startofpacket;                                                                // rsp_xbar_demux:src3_startofpacket -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_demux_src3_data;                                                                         // rsp_xbar_demux:src3_data -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] rsp_xbar_demux_src3_channel;                                                                      // rsp_xbar_demux:src3_channel -> 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src4_endofpacket;                                                                  // rsp_xbar_demux:src4_endofpacket -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src4_valid;                                                                        // rsp_xbar_demux:src4_valid -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src4_startofpacket;                                                                // rsp_xbar_demux:src4_startofpacket -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_demux_src4_data;                                                                         // rsp_xbar_demux:src4_data -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] rsp_xbar_demux_src4_channel;                                                                      // rsp_xbar_demux:src4_channel -> buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                            // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [83:0] addr_router_src_data;                                                                             // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [4:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_demux_src0_ready;                                                                        // p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire         addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [83:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [4:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_demux_src1_ready;                                                                        // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src1_ready
	wire         addr_router_002_src_endofpacket;                                                                  // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         addr_router_002_src_valid;                                                                        // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire         addr_router_002_src_startofpacket;                                                                // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [83:0] addr_router_002_src_data;                                                                         // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [4:0] addr_router_002_src_channel;                                                                      // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire         addr_router_002_src_ready;                                                                        // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire         rsp_xbar_demux_src2_ready;                                                                        // 3Dlizer_avalon_master_w_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src2_ready
	wire         addr_router_003_src_endofpacket;                                                                  // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         addr_router_003_src_valid;                                                                        // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire         addr_router_003_src_startofpacket;                                                                // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [83:0] addr_router_003_src_data;                                                                         // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [4:0] addr_router_003_src_channel;                                                                      // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire         addr_router_003_src_ready;                                                                        // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire         rsp_xbar_demux_src3_ready;                                                                        // 3Dlizer_avalon_master_r_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src3_ready
	wire         addr_router_004_src_endofpacket;                                                                  // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire         addr_router_004_src_valid;                                                                        // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire         addr_router_004_src_startofpacket;                                                                // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [83:0] addr_router_004_src_data;                                                                         // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [4:0] addr_router_004_src_channel;                                                                      // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire         addr_router_004_src_ready;                                                                        // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire         rsp_xbar_demux_src4_ready;                                                                        // buffer_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src4_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                           // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [83:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [4:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready

	nios_system_clocks clocks (
		.CLOCK_50    (clock_50_clk),                   //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),             //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.VGA_CLK     (clocks_vga_clk_clk)              //              vga_clk.clk
	);

	nios_system_v_decoder v_decoder (
		.clk                      (clocks_sys_clk_clk),                            //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),            //     clock_reset_reset.reset
		.stream_out_ready         (v_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (v_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (v_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (v_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (v_decoder_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_decoder_TD_CLK27),                        //    external_interface.export
		.TD_DATA                  (video_decoder_TD_DATA),                         //                      .export
		.TD_HS                    (video_decoder_TD_HS),                           //                      .export
		.TD_VS                    (video_decoder_TD_VS),                           //                      .export
		.clk27_reset              (video_decoder_clk27_reset),                     //                      .export
		.TD_RESET                 (video_decoder_TD_RESET),                        //                      .export
		.overflow_flag            (video_decoder_overflow_flag)                    //                      .export
	);

	nios_system_chroma_resampler chroma_resampler (
		.clk                      (clocks_sys_clk_clk),                                  //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                  //    clock_reset_reset.reset
		.stream_in_startofpacket  (v_decoder_avalon_decoder_source_startofpacket),       //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (v_decoder_avalon_decoder_source_endofpacket),         //                     .endofpacket
		.stream_in_valid          (v_decoder_avalon_decoder_source_valid),               //                     .valid
		.stream_in_ready          (v_decoder_avalon_decoder_source_ready),               //                     .ready
		.stream_in_data           (v_decoder_avalon_decoder_source_data),                //                     .data
		.stream_out_ready         (chroma_resampler_avalon_chroma_source_ready),         // avalon_chroma_source.ready
		.stream_out_startofpacket (chroma_resampler_avalon_chroma_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (chroma_resampler_avalon_chroma_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (chroma_resampler_avalon_chroma_source_valid),         //                     .valid
		.stream_out_data          (chroma_resampler_avalon_chroma_source_data)           //                     .data
	);

	nios_system_color_space_converter color_space_converter (
		.clk                      (clocks_sys_clk_clk),                                    //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                    // clock_reset_reset.reset
		.stream_in_startofpacket  (chroma_resampler_avalon_chroma_source_startofpacket),   //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (chroma_resampler_avalon_chroma_source_endofpacket),     //                  .endofpacket
		.stream_in_valid          (chroma_resampler_avalon_chroma_source_valid),           //                  .valid
		.stream_in_ready          (chroma_resampler_avalon_chroma_source_ready),           //                  .ready
		.stream_in_data           (chroma_resampler_avalon_chroma_source_data),            //                  .data
		.stream_out_ready         (color_space_converter_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (color_space_converter_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (color_space_converter_avalon_csc_source_data)           //                  .data
	);

	nios_system_v_rgb_resampler v_rgb_resampler (
		.clk                      (clocks_sys_clk_clk),                                    //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                    // clock_reset_reset.reset
		.stream_in_startofpacket  (color_space_converter_avalon_csc_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_in_ready          (color_space_converter_avalon_csc_source_ready),         //                  .ready
		.stream_in_data           (color_space_converter_avalon_csc_source_data),          //                  .data
		.stream_out_ready         (v_rgb_resampler_avalon_rgb_source_ready),               // avalon_rgb_source.ready
		.stream_out_startofpacket (v_rgb_resampler_avalon_rgb_source_startofpacket),       //                  .startofpacket
		.stream_out_endofpacket   (v_rgb_resampler_avalon_rgb_source_endofpacket),         //                  .endofpacket
		.stream_out_valid         (v_rgb_resampler_avalon_rgb_source_valid),               //                  .valid
		.stream_out_data          (v_rgb_resampler_avalon_rgb_source_data)                 //                  .data
	);

	nios_system_v_clipper v_clipper (
		.clk                      (clocks_sys_clk_clk),                              //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              //     clock_reset_reset.reset
		.stream_in_data           (v_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (v_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (v_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (v_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (v_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (v_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (v_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (v_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (v_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (v_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	nios_system_v_scaler v_scaler (
		.clk                      (clocks_sys_clk_clk),                            //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),            //    clock_reset_reset.reset
		.stream_in_startofpacket  (v_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (v_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (v_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (v_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (v_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (v_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (v_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (v_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (v_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (v_scaler_avalon_scaler_source_data)             //                     .data
	);

	nios_system_v_dma_controller v_dma_controller (
		.clk                  (clocks_sys_clk_clk),                             //              clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),             //        clock_reset_reset.reset
		.stream_data          (v_scaler_avalon_scaler_source_data),             //          avalon_dma_sink.data
		.stream_startofpacket (v_scaler_avalon_scaler_source_startofpacket),    //                         .startofpacket
		.stream_endofpacket   (v_scaler_avalon_scaler_source_endofpacket),      //                         .endofpacket
		.stream_valid         (v_scaler_avalon_scaler_source_valid),            //                         .valid
		.stream_ready         (v_scaler_avalon_scaler_source_ready),            //                         .ready
		.slave_address        (),                                               // avalon_dma_control_slave.address
		.slave_byteenable     (),                                               //                         .byteenable
		.slave_read           (),                                               //                         .read
		.slave_write          (),                                               //                         .write
		.slave_writedata      (),                                               //                         .writedata
		.slave_readdata       (),                                               //                         .readdata
		.master_address       (v_dma_controller_avalon_dma_master_address),     //        avalon_dma_master.address
		.master_waitrequest   (v_dma_controller_avalon_dma_master_waitrequest), //                         .waitrequest
		.master_write         (v_dma_controller_avalon_dma_master_write),       //                         .write
		.master_writedata     (v_dma_controller_avalon_dma_master_writedata)    //                         .writedata
	);

	nios_system_p_buffer_dma p_buffer_dma (
		.clk                  (clocks_sys_clk_clk),                                 //             clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),                 //       clock_reset_reset.reset
		.master_readdatavalid (p_buffer_dma_avalon_pixel_dma_master_readdatavalid), // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (p_buffer_dma_avalon_pixel_dma_master_waitrequest),   //                        .waitrequest
		.master_address       (p_buffer_dma_avalon_pixel_dma_master_address),       //                        .address
		.master_arbiterlock   (p_buffer_dma_avalon_pixel_dma_master_lock),          //                        .lock
		.master_read          (p_buffer_dma_avalon_pixel_dma_master_read),          //                        .read
		.master_readdata      (p_buffer_dma_avalon_pixel_dma_master_readdata),      //                        .readdata
		.slave_address        (),                                                   //    avalon_control_slave.address
		.slave_byteenable     (),                                                   //                        .byteenable
		.slave_read           (),                                                   //                        .read
		.slave_write          (),                                                   //                        .write
		.slave_writedata      (),                                                   //                        .writedata
		.slave_readdata       (),                                                   //                        .readdata
		.stream_ready         (p_buffer_dma_avalon_pixel_source_ready),             //     avalon_pixel_source.ready
		.stream_startofpacket (p_buffer_dma_avalon_pixel_source_startofpacket),     //                        .startofpacket
		.stream_endofpacket   (p_buffer_dma_avalon_pixel_source_endofpacket),       //                        .endofpacket
		.stream_valid         (p_buffer_dma_avalon_pixel_source_valid),             //                        .valid
		.stream_data          (p_buffer_dma_avalon_pixel_source_data)               //                        .data
	);

	nios_system_p_rgb_resampler p_rgb_resampler (
		.clk                      (clocks_sys_clk_clk),                              //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              // clock_reset_reset.reset
		.stream_in_startofpacket  (p_buffer_dma_avalon_pixel_source_startofpacket),  //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (p_buffer_dma_avalon_pixel_source_endofpacket),    //                  .endofpacket
		.stream_in_valid          (p_buffer_dma_avalon_pixel_source_valid),          //                  .valid
		.stream_in_ready          (p_buffer_dma_avalon_pixel_source_ready),          //                  .ready
		.stream_in_data           (p_buffer_dma_avalon_pixel_source_data),           //                  .data
		.stream_out_ready         (p_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (p_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (p_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (p_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (p_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_p_scaler p_scaler (
		.clk                      (clocks_sys_clk_clk),                              //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              //    clock_reset_reset.reset
		.stream_in_startofpacket  (p_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (p_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (p_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (p_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (p_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (p_scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (p_scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (p_scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (p_scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (p_scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_dual_clock_fifo dual_clock_fifo (
		.clk_stream_in            (clocks_sys_clk_clk),                                    //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                    //   clock_stream_in_reset.reset
		.clk_stream_out           (clocks_vga_clk_clk),                                    //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                    //  clock_stream_out_reset.reset
		.stream_in_ready          (p_scaler_avalon_scaler_source_ready),                   //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (p_scaler_avalon_scaler_source_startofpacket),           //                        .startofpacket
		.stream_in_endofpacket    (p_scaler_avalon_scaler_source_endofpacket),             //                        .endofpacket
		.stream_in_valid          (p_scaler_avalon_scaler_source_valid),                   //                        .valid
		.stream_in_data           (p_scaler_avalon_scaler_source_data),                    //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_vga_controller vga_controller (
		.clk           (clocks_vga_clk_clk),                                    //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),                    //  clock_reset_reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                                    // external_interface.export
		.VGA_HS        (vga_controller_HS),                                     //                   .export
		.VGA_VS        (vga_controller_VS),                                     //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                                  //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                                   //                   .export
		.VGA_R         (vga_controller_R),                                      //                   .export
		.VGA_G         (vga_controller_G),                                      //                   .export
		.VGA_B         (vga_controller_B)                                       //                   .export
	);

	nios_system_p_buffer p_buffer (
		.clk           (clocks_sys_clk_clk),                                                      //        clock_reset.clk
		.reset         (rst_controller_001_reset_out_reset),                                      //  clock_reset_reset.reset
		.SRAM_DQ       (sram_DQ),                                                                 // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                               //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                               //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                               //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                               //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                               //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                               //                   .export
		.address       (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	threeDlizer #(
		.pixel_buffer_2D (32'b00000000000000000000000000000000),
		.pixel_buffer_3D (32'b00000000000000100101100000000000)
	) id3dlizer (
		.reset_out     (threedlizer_reset_out),                 //     conduit_end.export
		.pixel_r_ready (threedlizer_pixel_r_ready),             //                .export
		.pixel_r       (threedlizer_pixel_r),                   //                .export
		.pixel_offset  (threedlizer_pixel_offset),              //                .export
		.pixel_r_done  (threedlizer_pixel_r_done),              //                .export
		.red_led       (threedlizer_red_led),                   //                .export
		.clk_in        (threedlizer_clk_in),                    //                .export
		.clk           (clocks_sys_clk_clk),                    //           clock.clk
		.reset_in      (~rst_controller_001_reset_out_reset),   //           reset.reset_n
		.master_wr_en  (id3dlizer_avalon_master_w_write),       // avalon_master_w.write
		.master_wd     (id3dlizer_avalon_master_w_writedata),   //                .writedata
		.master_w_wait (id3dlizer_avalon_master_w_waitrequest), //                .waitrequest
		.master_w_addr (id3dlizer_avalon_master_w_address),     //                .address
		.master_w_be   (id3dlizer_avalon_master_w_byteenable),  //                .byteenable
		.master_rd     (id3dlizer_avalon_master_r_readdata),    // avalon_master_r.readdata
		.master_rd_en  (id3dlizer_avalon_master_r_read),        //                .read
		.master_r_wait (id3dlizer_avalon_master_r_waitrequest), //                .waitrequest
		.master_r_addr (id3dlizer_avalon_master_r_address),     //                .address
		.master_r_be   (id3dlizer_avalon_master_r_byteenable)   //                .byteenable
	);

	buffer_reader #(
		.pixel_buffer_base (32'b00000000000000100101100000000000)
	) buffer_reader (
		.clk           (clocks_sys_clk_clk),                      //         clock.clk
		.clk_in        (buffer_reader_clk_in),                    //   conduit_end.export
		.pixel_set     (buffer_reader_pixel_set),                 //              .export
		.pixel_offset  (buffer_reader_pixel_offset),              //              .export
		.pixel_ready   (buffer_reader_pixel_ready),               //              .export
		.pixel         (buffer_reader_pixel),                     //              .export
		.red_led       (buffer_reader_red_led),                   //              .export
		.master_r_wait (buffer_reader_avalon_master_waitrequest), // avalon_master.waitrequest
		.master_rd_en  (buffer_reader_avalon_master_read),        //              .read
		.master_rd     (buffer_reader_avalon_master_readdata),    //              .readdata
		.master_r_addr (buffer_reader_avalon_master_address),     //              .address
		.master_r_be   (buffer_reader_avalon_master_byteenable),  //              .byteenable
		.rst           (~rst_controller_001_reset_out_reset)      //         reset.reset_n
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) p_buffer_dma_avalon_pixel_dma_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                      //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                      //                     reset.reset
		.uav_address              (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (p_buffer_dma_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (p_buffer_dma_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (p_buffer_dma_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata              (p_buffer_dma_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (p_buffer_dma_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (p_buffer_dma_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                    //               (terminated)
		.av_byteenable            (2'b11),                                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                                    //               (terminated)
		.av_write                 (1'b0),                                                                                    //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                                    //               (terminated)
		.uav_clken                (),                                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                                   //               (terminated)
		.av_response              (),                                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) v_dma_controller_avalon_dma_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                     reset.reset
		.uav_address              (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (v_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (v_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write                 (v_dma_controller_avalon_dma_master_write),                                              //                          .write
		.av_writedata             (v_dma_controller_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                  //               (terminated)
		.av_byteenable            (2'b11),                                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                                  //               (terminated)
		.av_read                  (1'b0),                                                                                  //               (terminated)
		.av_readdata              (),                                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                                  //               (terminated)
		.uav_clken                (),                                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                                 //               (terminated)
		.av_response              (),                                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) id3dlizer_avalon_master_w_translator (
		.clk                      (clocks_sys_clk_clk),                                                           //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address              (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (id3dlizer_avalon_master_w_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (id3dlizer_avalon_master_w_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (id3dlizer_avalon_master_w_byteenable),                                         //                          .byteenable
		.av_write                 (id3dlizer_avalon_master_w_write),                                              //                          .write
		.av_writedata             (id3dlizer_avalon_master_w_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                         //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_read                  (1'b0),                                                                         //               (terminated)
		.av_readdata              (),                                                                             //               (terminated)
		.av_readdatavalid         (),                                                                             //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.av_debugaccess           (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) id3dlizer_avalon_master_r_translator (
		.clk                      (clocks_sys_clk_clk),                                                           //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address              (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (id3dlizer_avalon_master_r_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (id3dlizer_avalon_master_r_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (id3dlizer_avalon_master_r_byteenable),                                         //                          .byteenable
		.av_read                  (id3dlizer_avalon_master_r_read),                                               //                          .read
		.av_readdata              (id3dlizer_avalon_master_r_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                         //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_readdatavalid         (),                                                                             //               (terminated)
		.av_write                 (1'b0),                                                                         //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                         //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.av_debugaccess           (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) buffer_reader_avalon_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                     reset.reset
		.uav_address              (buffer_reader_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (buffer_reader_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (buffer_reader_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (buffer_reader_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (buffer_reader_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (buffer_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (buffer_reader_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (buffer_reader_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (buffer_reader_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (buffer_reader_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (buffer_reader_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (buffer_reader_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (buffer_reader_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (buffer_reader_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (buffer_reader_avalon_master_read),                                               //                          .read
		.av_readdata              (buffer_reader_avalon_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) p_buffer_avalon_sram_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.av_address              (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src0_valid),                                                                        //        rp.valid
		.rp_data                 (rsp_xbar_demux_src0_data),                                                                         //          .data
		.rp_channel              (rsp_xbar_demux_src0_channel),                                                                      //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src0_startofpacket),                                                                //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src0_endofpacket),                                                                  //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src0_ready),                                                                        //          .ready
		.av_response             (),                                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.av_address              (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src1_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_demux_src1_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_demux_src1_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src1_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src1_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src1_ready),                                                                      //          .ready
		.av_response             (),                                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address              (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src2_valid),                                                             //        rp.valid
		.rp_data                 (rsp_xbar_demux_src2_data),                                                              //          .data
		.rp_channel              (rsp_xbar_demux_src2_channel),                                                           //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src2_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src2_endofpacket),                                                       //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src2_ready),                                                             //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address              (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src3_valid),                                                             //        rp.valid
		.rp_data                 (rsp_xbar_demux_src3_data),                                                              //          .data
		.rp_channel              (rsp_xbar_demux_src3_channel),                                                           //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src3_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src3_endofpacket),                                                       //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src3_ready),                                                             //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_THREAD_ID_H           (74),
		.PKT_THREAD_ID_L           (74),
		.PKT_CACHE_H               (81),
		.PKT_CACHE_L               (78),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) buffer_reader_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.av_address              (buffer_reader_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (buffer_reader_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (buffer_reader_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (buffer_reader_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (buffer_reader_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (buffer_reader_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (buffer_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (buffer_reader_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (buffer_reader_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (buffer_reader_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (buffer_reader_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src4_valid),                                                               //        rp.valid
		.rp_data                 (rsp_xbar_demux_src4_data),                                                                //          .data
		.rp_channel              (rsp_xbar_demux_src4_channel),                                                             //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src4_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src4_endofpacket),                                                         //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src4_ready),                                                               //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                        //                .channel
		.rf_sink_ready           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (p_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                            //       src.ready
		.src_valid          (addr_router_src_valid),                                                                            //          .valid
		.src_data           (addr_router_src_data),                                                                             //          .data
		.src_channel        (addr_router_src_channel),                                                                          //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                       //          .endofpacket
	);

	nios_system_addr_router addr_router_001 (
		.sink_ready         (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                      //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                      //          .valid
		.src_data           (addr_router_001_src_data),                                                                       //          .data
		.src_channel        (addr_router_001_src_channel),                                                                    //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_system_addr_router addr_router_002 (
		.sink_ready         (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (id3dlizer_avalon_master_w_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                             //          .valid
		.src_data           (addr_router_002_src_data),                                                              //          .data
		.src_channel        (addr_router_002_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_addr_router addr_router_003 (
		.sink_ready         (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (id3dlizer_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_addr_router addr_router_004 (
		.sink_ready         (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (buffer_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                               //          .valid
		.src_data           (addr_router_004_src_data),                                                                //          .data
		.src_channel        (addr_router_004_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_50_reset_n),              // reset_in0.reset
		.clk        (clock_50_clk),                   //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_50_reset_n),                  // reset_in0.reset
		.clk        (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_50_reset_n),                  // reset_in0.reset
		.clk        (clocks_vga_clk_clk),                 //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready         (rsp_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid         (rsp_xbar_demux_src2_valid),          //          .valid
		.src2_data          (rsp_xbar_demux_src2_data),           //          .data
		.src2_channel       (rsp_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket (rsp_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready         (rsp_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid         (rsp_xbar_demux_src3_valid),          //          .valid
		.src3_data          (rsp_xbar_demux_src3_data),           //          .data
		.src3_channel       (rsp_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket (rsp_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_src3_endofpacket),    //          .endofpacket
		.src4_ready         (rsp_xbar_demux_src4_ready),          //      src4.ready
		.src4_valid         (rsp_xbar_demux_src4_valid),          //          .valid
		.src4_data          (rsp_xbar_demux_src4_data),           //          .data
		.src4_channel       (rsp_xbar_demux_src4_channel),        //          .channel
		.src4_startofpacket (rsp_xbar_demux_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_src4_endofpacket)     //          .endofpacket
	);

endmodule
