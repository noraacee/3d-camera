// nios_system.v

// Generated using ACDS version 13.0sp1 232 at 2015.04.08.19:36:37

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clock_50_clk,                //      clock_50.clk
		input  wire        reset_50_reset_n,            //      reset_50.reset_n
		input  wire        video_decoder_TD_CLK27,      // video_decoder.TD_CLK27
		input  wire [7:0]  video_decoder_TD_DATA,       //              .TD_DATA
		input  wire        video_decoder_TD_HS,         //              .TD_HS
		input  wire        video_decoder_TD_VS,         //              .TD_VS
		input  wire        video_decoder_clk27_reset,   //              .clk27_reset
		output wire        video_decoder_TD_RESET,      //              .TD_RESET
		output wire        video_decoder_overflow_flag, //              .overflow_flag
		inout  wire [15:0] sram_DQ,                     //          sram.DQ
		output wire [17:0] sram_ADDR,                   //              .ADDR
		output wire        sram_LB_N,                   //              .LB_N
		output wire        sram_UB_N,                   //              .UB_N
		output wire        sram_CE_N,                   //              .CE_N
		output wire        sram_OE_N,                   //              .OE_N
		output wire        sram_WE_N,                   //              .WE_N
		output wire        red_extractor_pixel_r_ready, // red_extractor.pixel_r_ready
		output wire [4:0]  red_extractor_pixel_r,       //              .pixel_r
		output wire [17:0] red_extractor_pixel_offset,  //              .pixel_offset
		input  wire        red_extractor_reset_in,      //              .reset_in
		output wire [17:0] red_extractor_red_led,       //              .red_led
		input  wire        red_extractor_pixel_r_done,  //              .pixel_r_done
		input  wire        red_extractor_clk_in         //              .clk_in
	);

	wire         clocks_sys_clk_clk;                                                                              // clocks:sys_clk -> [addr_router:clk, addr_router_001:clk, chroma_resampler:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, color_space_converter:clk, id_router:clk, p_buffer:clk, p_buffer_avalon_sram_slave_translator:clk, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, red_extractor:clk, red_extractor_avalon_master_r_translator:clk, red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux:clk, rst_controller_001:clk, v_clipper:clk, v_decoder:clk, v_dma_controller:clk, v_dma_controller_avalon_dma_master_translator:clk, v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, v_rgb_resampler:clk, v_scaler:clk]
	wire         v_decoder_avalon_decoder_source_endofpacket;                                                     // v_decoder:stream_out_endofpacket -> chroma_resampler:stream_in_endofpacket
	wire         v_decoder_avalon_decoder_source_valid;                                                           // v_decoder:stream_out_valid -> chroma_resampler:stream_in_valid
	wire         v_decoder_avalon_decoder_source_startofpacket;                                                   // v_decoder:stream_out_startofpacket -> chroma_resampler:stream_in_startofpacket
	wire  [15:0] v_decoder_avalon_decoder_source_data;                                                            // v_decoder:stream_out_data -> chroma_resampler:stream_in_data
	wire         v_decoder_avalon_decoder_source_ready;                                                           // chroma_resampler:stream_in_ready -> v_decoder:stream_out_ready
	wire         chroma_resampler_avalon_chroma_source_endofpacket;                                               // chroma_resampler:stream_out_endofpacket -> color_space_converter:stream_in_endofpacket
	wire         chroma_resampler_avalon_chroma_source_valid;                                                     // chroma_resampler:stream_out_valid -> color_space_converter:stream_in_valid
	wire         chroma_resampler_avalon_chroma_source_startofpacket;                                             // chroma_resampler:stream_out_startofpacket -> color_space_converter:stream_in_startofpacket
	wire  [23:0] chroma_resampler_avalon_chroma_source_data;                                                      // chroma_resampler:stream_out_data -> color_space_converter:stream_in_data
	wire         chroma_resampler_avalon_chroma_source_ready;                                                     // color_space_converter:stream_in_ready -> chroma_resampler:stream_out_ready
	wire         color_space_converter_avalon_csc_source_endofpacket;                                             // color_space_converter:stream_out_endofpacket -> v_rgb_resampler:stream_in_endofpacket
	wire         color_space_converter_avalon_csc_source_valid;                                                   // color_space_converter:stream_out_valid -> v_rgb_resampler:stream_in_valid
	wire         color_space_converter_avalon_csc_source_startofpacket;                                           // color_space_converter:stream_out_startofpacket -> v_rgb_resampler:stream_in_startofpacket
	wire  [23:0] color_space_converter_avalon_csc_source_data;                                                    // color_space_converter:stream_out_data -> v_rgb_resampler:stream_in_data
	wire         color_space_converter_avalon_csc_source_ready;                                                   // v_rgb_resampler:stream_in_ready -> color_space_converter:stream_out_ready
	wire         v_rgb_resampler_avalon_rgb_source_endofpacket;                                                   // v_rgb_resampler:stream_out_endofpacket -> v_clipper:stream_in_endofpacket
	wire         v_rgb_resampler_avalon_rgb_source_valid;                                                         // v_rgb_resampler:stream_out_valid -> v_clipper:stream_in_valid
	wire         v_rgb_resampler_avalon_rgb_source_startofpacket;                                                 // v_rgb_resampler:stream_out_startofpacket -> v_clipper:stream_in_startofpacket
	wire  [15:0] v_rgb_resampler_avalon_rgb_source_data;                                                          // v_rgb_resampler:stream_out_data -> v_clipper:stream_in_data
	wire         v_rgb_resampler_avalon_rgb_source_ready;                                                         // v_clipper:stream_in_ready -> v_rgb_resampler:stream_out_ready
	wire         v_clipper_avalon_clipper_source_endofpacket;                                                     // v_clipper:stream_out_endofpacket -> v_scaler:stream_in_endofpacket
	wire         v_clipper_avalon_clipper_source_valid;                                                           // v_clipper:stream_out_valid -> v_scaler:stream_in_valid
	wire         v_clipper_avalon_clipper_source_startofpacket;                                                   // v_clipper:stream_out_startofpacket -> v_scaler:stream_in_startofpacket
	wire  [15:0] v_clipper_avalon_clipper_source_data;                                                            // v_clipper:stream_out_data -> v_scaler:stream_in_data
	wire         v_clipper_avalon_clipper_source_ready;                                                           // v_scaler:stream_in_ready -> v_clipper:stream_out_ready
	wire         v_scaler_avalon_scaler_source_endofpacket;                                                       // v_scaler:stream_out_endofpacket -> v_dma_controller:stream_endofpacket
	wire         v_scaler_avalon_scaler_source_valid;                                                             // v_scaler:stream_out_valid -> v_dma_controller:stream_valid
	wire         v_scaler_avalon_scaler_source_startofpacket;                                                     // v_scaler:stream_out_startofpacket -> v_dma_controller:stream_startofpacket
	wire  [15:0] v_scaler_avalon_scaler_source_data;                                                              // v_scaler:stream_out_data -> v_dma_controller:stream_data
	wire         v_scaler_avalon_scaler_source_ready;                                                             // v_dma_controller:stream_ready -> v_scaler:stream_out_ready
	wire         v_dma_controller_avalon_dma_master_waitrequest;                                                  // v_dma_controller_avalon_dma_master_translator:av_waitrequest -> v_dma_controller:master_waitrequest
	wire  [15:0] v_dma_controller_avalon_dma_master_writedata;                                                    // v_dma_controller:master_writedata -> v_dma_controller_avalon_dma_master_translator:av_writedata
	wire  [31:0] v_dma_controller_avalon_dma_master_address;                                                      // v_dma_controller:master_address -> v_dma_controller_avalon_dma_master_translator:av_address
	wire         v_dma_controller_avalon_dma_master_write;                                                        // v_dma_controller:master_write -> v_dma_controller_avalon_dma_master_translator:av_write
	wire         red_extractor_avalon_master_r_waitrequest;                                                       // red_extractor_avalon_master_r_translator:av_waitrequest -> red_extractor:master_r_wait
	wire  [31:0] red_extractor_avalon_master_r_address;                                                           // red_extractor:master_r_addr -> red_extractor_avalon_master_r_translator:av_address
	wire         red_extractor_avalon_master_r_read;                                                              // red_extractor:master_rd_en -> red_extractor_avalon_master_r_translator:av_read
	wire  [15:0] red_extractor_avalon_master_r_readdata;                                                          // red_extractor_avalon_master_r_translator:av_readdata -> red_extractor:master_rd
	wire   [1:0] red_extractor_avalon_master_r_byteenable;                                                        // red_extractor:master_r_be -> red_extractor_avalon_master_r_translator:av_byteenable
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                             // p_buffer_avalon_sram_slave_translator:av_writedata -> p_buffer:writedata
	wire  [17:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                               // p_buffer_avalon_sram_slave_translator:av_address -> p_buffer:address
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                 // p_buffer_avalon_sram_slave_translator:av_write -> p_buffer:write
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                  // p_buffer_avalon_sram_slave_translator:av_read -> p_buffer:read
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                              // p_buffer:readdata -> p_buffer_avalon_sram_slave_translator:av_readdata
	wire         p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                         // p_buffer:readdatavalid -> p_buffer_avalon_sram_slave_translator:av_readdatavalid
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                            // p_buffer_avalon_sram_slave_translator:av_byteenable -> p_buffer:byteenable
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;             // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> v_dma_controller_avalon_dma_master_translator:uav_waitrequest
	wire   [1:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;              // v_dma_controller_avalon_dma_master_translator:uav_burstcount -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;               // v_dma_controller_avalon_dma_master_translator:uav_writedata -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                 // v_dma_controller_avalon_dma_master_translator:uav_address -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                    // v_dma_controller_avalon_dma_master_translator:uav_lock -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                   // v_dma_controller_avalon_dma_master_translator:uav_write -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                    // v_dma_controller_avalon_dma_master_translator:uav_read -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> v_dma_controller_avalon_dma_master_translator:uav_readdata
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;             // v_dma_controller_avalon_dma_master_translator:uav_debugaccess -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;              // v_dma_controller_avalon_dma_master_translator:uav_byteenable -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;           // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> v_dma_controller_avalon_dma_master_translator:uav_readdatavalid
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_waitrequest;                  // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_waitrequest -> red_extractor_avalon_master_r_translator:uav_waitrequest
	wire   [1:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_burstcount;                   // red_extractor_avalon_master_r_translator:uav_burstcount -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_writedata;                    // red_extractor_avalon_master_r_translator:uav_writedata -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_address;                      // red_extractor_avalon_master_r_translator:uav_address -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_address
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_lock;                         // red_extractor_avalon_master_r_translator:uav_lock -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_lock
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_write;                        // red_extractor_avalon_master_r_translator:uav_write -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_write
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_read;                         // red_extractor_avalon_master_r_translator:uav_read -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdata;                     // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_readdata -> red_extractor_avalon_master_r_translator:uav_readdata
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_debugaccess;                  // red_extractor_avalon_master_r_translator:uav_debugaccess -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_byteenable;                   // red_extractor_avalon_master_r_translator:uav_byteenable -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_byteenable
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdatavalid;                // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:av_readdatavalid -> red_extractor_avalon_master_r_translator:uav_readdatavalid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // p_buffer_avalon_sram_slave_translator:uav_waitrequest -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> p_buffer_avalon_sram_slave_translator:uav_burstcount
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> p_buffer_avalon_sram_slave_translator:uav_writedata
	wire  [31:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> p_buffer_avalon_sram_slave_translator:uav_address
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> p_buffer_avalon_sram_slave_translator:uav_write
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> p_buffer_avalon_sram_slave_translator:uav_lock
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> p_buffer_avalon_sram_slave_translator:uav_read
	wire  [15:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // p_buffer_avalon_sram_slave_translator:uav_readdata -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // p_buffer_avalon_sram_slave_translator:uav_readdatavalid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> p_buffer_avalon_sram_slave_translator:uav_debugaccess
	wire   [1:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> p_buffer_avalon_sram_slave_translator:uav_byteenable
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [80:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [80:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [17:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;    // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;          // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;  // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [79:0] v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;           // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;          // addr_router:sink_ready -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket;         // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid;               // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket;       // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [79:0] red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data;                // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready;               // addr_router_001:sink_ready -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:cp_ready
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [79:0] p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                  // rst_controller:reset_out -> clocks:reset
	wire         rst_controller_001_reset_out_reset;                                                              // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, chroma_resampler:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, color_space_converter:reset, id_router:reset, p_buffer:reset, p_buffer_avalon_sram_slave_translator:reset, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, red_extractor:reset_n_in, red_extractor_avalon_master_r_translator:reset, red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, v_clipper:reset, v_decoder:reset, v_dma_controller:reset, v_dma_controller_avalon_dma_master_translator:reset, v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, v_rgb_resampler:reset, v_scaler:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                 // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                       // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                               // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [79:0] cmd_xbar_demux_src0_data;                                                                        // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                     // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                       // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                             // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                   // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                           // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [79:0] cmd_xbar_demux_001_src0_data;                                                                    // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [1:0] cmd_xbar_demux_001_src0_channel;                                                                 // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                   // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                 // rsp_xbar_demux:src0_endofpacket -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                       // rsp_xbar_demux:src0_valid -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                               // rsp_xbar_demux:src0_startofpacket -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [79:0] rsp_xbar_demux_src0_data;                                                                        // rsp_xbar_demux:src0_data -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                     // rsp_xbar_demux:src0_channel -> v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src1_endofpacket;                                                                 // rsp_xbar_demux:src1_endofpacket -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                       // rsp_xbar_demux:src1_valid -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                               // rsp_xbar_demux:src1_startofpacket -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [79:0] rsp_xbar_demux_src1_data;                                                                        // rsp_xbar_demux:src1_data -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_src1_channel;                                                                     // rsp_xbar_demux:src1_channel -> red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_channel
	wire         addr_router_src_endofpacket;                                                                     // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                           // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                   // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [79:0] addr_router_src_data;                                                                            // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] addr_router_src_channel;                                                                         // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                           // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_demux_src0_ready;                                                                       // v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire         addr_router_001_src_endofpacket;                                                                 // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                       // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                               // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [79:0] addr_router_001_src_data;                                                                        // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [1:0] addr_router_001_src_channel;                                                                     // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                       // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_demux_src1_ready;                                                                       // red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src1_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                    // cmd_xbar_mux:src_endofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                          // cmd_xbar_mux:src_valid -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                  // cmd_xbar_mux:src_startofpacket -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [79:0] cmd_xbar_mux_src_data;                                                                           // cmd_xbar_mux:src_data -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_src_channel;                                                                        // cmd_xbar_mux:src_channel -> p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                          // p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                       // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                             // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                     // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [79:0] id_router_src_data;                                                                              // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                           // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                             // rsp_xbar_demux:sink_ready -> id_router:src_ready

	nios_system_clocks clocks (
		.CLOCK_50    (clock_50_clk),                   //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),             //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.VGA_CLK     ()                                //              vga_clk.clk
	);

	nios_system_v_decoder v_decoder (
		.clk                      (clocks_sys_clk_clk),                            //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),            //     clock_reset_reset.reset
		.stream_out_ready         (v_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (v_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (v_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (v_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (v_decoder_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_decoder_TD_CLK27),                        //    external_interface.export
		.TD_DATA                  (video_decoder_TD_DATA),                         //                      .export
		.TD_HS                    (video_decoder_TD_HS),                           //                      .export
		.TD_VS                    (video_decoder_TD_VS),                           //                      .export
		.clk27_reset              (video_decoder_clk27_reset),                     //                      .export
		.TD_RESET                 (video_decoder_TD_RESET),                        //                      .export
		.overflow_flag            (video_decoder_overflow_flag)                    //                      .export
	);

	nios_system_chroma_resampler chroma_resampler (
		.clk                      (clocks_sys_clk_clk),                                  //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                  //    clock_reset_reset.reset
		.stream_in_startofpacket  (v_decoder_avalon_decoder_source_startofpacket),       //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (v_decoder_avalon_decoder_source_endofpacket),         //                     .endofpacket
		.stream_in_valid          (v_decoder_avalon_decoder_source_valid),               //                     .valid
		.stream_in_ready          (v_decoder_avalon_decoder_source_ready),               //                     .ready
		.stream_in_data           (v_decoder_avalon_decoder_source_data),                //                     .data
		.stream_out_ready         (chroma_resampler_avalon_chroma_source_ready),         // avalon_chroma_source.ready
		.stream_out_startofpacket (chroma_resampler_avalon_chroma_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (chroma_resampler_avalon_chroma_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (chroma_resampler_avalon_chroma_source_valid),         //                     .valid
		.stream_out_data          (chroma_resampler_avalon_chroma_source_data)           //                     .data
	);

	nios_system_color_space_converter color_space_converter (
		.clk                      (clocks_sys_clk_clk),                                    //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                    // clock_reset_reset.reset
		.stream_in_startofpacket  (chroma_resampler_avalon_chroma_source_startofpacket),   //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (chroma_resampler_avalon_chroma_source_endofpacket),     //                  .endofpacket
		.stream_in_valid          (chroma_resampler_avalon_chroma_source_valid),           //                  .valid
		.stream_in_ready          (chroma_resampler_avalon_chroma_source_ready),           //                  .ready
		.stream_in_data           (chroma_resampler_avalon_chroma_source_data),            //                  .data
		.stream_out_ready         (color_space_converter_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (color_space_converter_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (color_space_converter_avalon_csc_source_data)           //                  .data
	);

	nios_system_v_rgb_resampler v_rgb_resampler (
		.clk                      (clocks_sys_clk_clk),                                    //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                    // clock_reset_reset.reset
		.stream_in_startofpacket  (color_space_converter_avalon_csc_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (color_space_converter_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (color_space_converter_avalon_csc_source_valid),         //                  .valid
		.stream_in_ready          (color_space_converter_avalon_csc_source_ready),         //                  .ready
		.stream_in_data           (color_space_converter_avalon_csc_source_data),          //                  .data
		.stream_out_ready         (v_rgb_resampler_avalon_rgb_source_ready),               // avalon_rgb_source.ready
		.stream_out_startofpacket (v_rgb_resampler_avalon_rgb_source_startofpacket),       //                  .startofpacket
		.stream_out_endofpacket   (v_rgb_resampler_avalon_rgb_source_endofpacket),         //                  .endofpacket
		.stream_out_valid         (v_rgb_resampler_avalon_rgb_source_valid),               //                  .valid
		.stream_out_data          (v_rgb_resampler_avalon_rgb_source_data)                 //                  .data
	);

	nios_system_v_clipper v_clipper (
		.clk                      (clocks_sys_clk_clk),                              //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              //     clock_reset_reset.reset
		.stream_in_data           (v_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (v_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (v_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (v_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (v_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (v_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (v_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (v_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (v_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (v_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	nios_system_v_scaler v_scaler (
		.clk                      (clocks_sys_clk_clk),                            //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),            //    clock_reset_reset.reset
		.stream_in_startofpacket  (v_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (v_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (v_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (v_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (v_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (v_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (v_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (v_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (v_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (v_scaler_avalon_scaler_source_data)             //                     .data
	);

	nios_system_v_dma_controller v_dma_controller (
		.clk                  (clocks_sys_clk_clk),                             //              clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),             //        clock_reset_reset.reset
		.stream_data          (v_scaler_avalon_scaler_source_data),             //          avalon_dma_sink.data
		.stream_startofpacket (v_scaler_avalon_scaler_source_startofpacket),    //                         .startofpacket
		.stream_endofpacket   (v_scaler_avalon_scaler_source_endofpacket),      //                         .endofpacket
		.stream_valid         (v_scaler_avalon_scaler_source_valid),            //                         .valid
		.stream_ready         (v_scaler_avalon_scaler_source_ready),            //                         .ready
		.slave_address        (),                                               // avalon_dma_control_slave.address
		.slave_byteenable     (),                                               //                         .byteenable
		.slave_read           (),                                               //                         .read
		.slave_write          (),                                               //                         .write
		.slave_writedata      (),                                               //                         .writedata
		.slave_readdata       (),                                               //                         .readdata
		.master_address       (v_dma_controller_avalon_dma_master_address),     //        avalon_dma_master.address
		.master_waitrequest   (v_dma_controller_avalon_dma_master_waitrequest), //                         .waitrequest
		.master_write         (v_dma_controller_avalon_dma_master_write),       //                         .write
		.master_writedata     (v_dma_controller_avalon_dma_master_writedata)    //                         .writedata
	);

	nios_system_p_buffer p_buffer (
		.clk           (clocks_sys_clk_clk),                                                      //        clock_reset.clk
		.reset         (rst_controller_001_reset_out_reset),                                      //  clock_reset_reset.reset
		.SRAM_DQ       (sram_DQ),                                                                 // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                               //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                               //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                               //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                               //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                               //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                               //                   .export
		.address       (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	red_extractor #(
		.pixel_buffer_base (32'b00000000000000000000000000000000)
	) red_extractor (
		.clk           (clocks_sys_clk_clk),                        //           clock.clk
		.pixel_r_ready (red_extractor_pixel_r_ready),               //     conduit_end.export
		.pixel_r       (red_extractor_pixel_r),                     //                .export
		.pixel_offset  (red_extractor_pixel_offset),                //                .export
		.reset_in      (red_extractor_reset_in),                    //                .export
		.red_led       (red_extractor_red_led),                     //                .export
		.pixel_r_done  (red_extractor_pixel_r_done),                //                .export
		.clk_in        (red_extractor_clk_in),                      //                .export
		.reset_n_in    (~rst_controller_001_reset_out_reset),       //           reset.reset_n
		.master_rd     (red_extractor_avalon_master_r_readdata),    // avalon_master_r.readdata
		.master_rd_en  (red_extractor_avalon_master_r_read),        //                .read
		.master_r_wait (red_extractor_avalon_master_r_waitrequest), //                .waitrequest
		.master_r_addr (red_extractor_avalon_master_r_address),     //                .address
		.master_r_be   (red_extractor_avalon_master_r_byteenable)   //                .byteenable
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) v_dma_controller_avalon_dma_master_translator (
		.clk                      (clocks_sys_clk_clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                     reset.reset
		.uav_address              (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (v_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (v_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write                 (v_dma_controller_avalon_dma_master_write),                                              //                          .write
		.av_writedata             (v_dma_controller_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                  //               (terminated)
		.av_byteenable            (2'b11),                                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                                  //               (terminated)
		.av_read                  (1'b0),                                                                                  //               (terminated)
		.av_readdata              (),                                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                                  //               (terminated)
		.uav_clken                (),                                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                                 //               (terminated)
		.av_response              (),                                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) red_extractor_avalon_master_r_translator (
		.clk                      (clocks_sys_clk_clk),                                                               //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                               //                     reset.reset
		.uav_address              (red_extractor_avalon_master_r_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (red_extractor_avalon_master_r_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (red_extractor_avalon_master_r_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (red_extractor_avalon_master_r_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (red_extractor_avalon_master_r_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (red_extractor_avalon_master_r_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (red_extractor_avalon_master_r_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (red_extractor_avalon_master_r_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (red_extractor_avalon_master_r_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (red_extractor_avalon_master_r_byteenable),                                         //                          .byteenable
		.av_read                  (red_extractor_avalon_master_r_read),                                               //                          .read
		.av_readdata              (red_extractor_avalon_master_r_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_readdatavalid         (),                                                                                 //               (terminated)
		.av_write                 (1'b0),                                                                             //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) p_buffer_avalon_sram_slave_translator (
		.clk                      (clocks_sys_clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (p_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (70),
		.PKT_THREAD_ID_L           (70),
		.PKT_CACHE_H               (77),
		.PKT_CACHE_L               (74),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.av_address              (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src0_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_demux_src0_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_demux_src0_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src0_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src0_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src0_ready),                                                                      //          .ready
		.av_response             (),                                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (70),
		.PKT_THREAD_ID_L           (70),
		.PKT_CACHE_H               (77),
		.PKT_CACHE_L               (74),
		.PKT_DATA_SIDEBAND_H       (65),
		.PKT_DATA_SIDEBAND_L       (65),
		.PKT_QOS_H                 (67),
		.PKT_QOS_L                 (67),
		.PKT_ADDR_SIDEBAND_H       (64),
		.PKT_ADDR_SIDEBAND_L       (64),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.av_address              (red_extractor_avalon_master_r_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (red_extractor_avalon_master_r_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (red_extractor_avalon_master_r_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (red_extractor_avalon_master_r_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (red_extractor_avalon_master_r_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (red_extractor_avalon_master_r_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (red_extractor_avalon_master_r_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (red_extractor_avalon_master_r_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src1_valid),                                                                 //        rp.valid
		.rp_data                 (rsp_xbar_demux_src1_data),                                                                  //          .data
		.rp_channel              (rsp_xbar_demux_src1_channel),                                                               //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src1_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src1_endofpacket),                                                           //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src1_ready),                                                                 //          .ready
		.av_response             (),                                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                        //                .channel
		.rf_sink_ready           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (v_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                                          //          .valid
		.src_data           (addr_router_src_data),                                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_addr_router addr_router_001 (
		.sink_ready         (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (red_extractor_avalon_master_r_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                 //          .valid
		.src_data           (addr_router_001_src_data),                                                                  //          .data
		.src_channel        (addr_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (p_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_50_reset_n),              // reset_in0.reset
		.clk        (clock_50_clk),                   //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_50_reset_n),                  // reset_in0.reset
		.clk        (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

endmodule
